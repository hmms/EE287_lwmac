module lwmac(clk,reset,busWrite,busDataToLmac,busDataFromLmac,busAddr,pushSym,Sym,pushOut,dataOut,macSate);
input

endmodule